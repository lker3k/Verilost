
module vga (
	clk_clk,
	filter_mode_filter_mode,
	reset_reset_n,
	vga_CLK,
	vga_HS,
	vga_VS,
	vga_BLANK,
	vga_SYNC,
	vga_R,
	vga_G,
	vga_B,
	x_ready_x_ready);	

	input		clk_clk;
	input	[2:0]	filter_mode_filter_mode;
	input		reset_reset_n;
	output		vga_CLK;
	output		vga_HS;
	output		vga_VS;
	output		vga_BLANK;
	output		vga_SYNC;
	output	[7:0]	vga_R;
	output	[7:0]	vga_G;
	output	[7:0]	vga_B;
	output		x_ready_x_ready;
endmodule
